`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:23:09 08/03/2017 
// Design Name: 
// Module Name:    readoutSM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module readoutSM(
    output reg [7:0] ROWADD,  //see timing diagram for signal definitions
    output reg COL_L_EN,
    output reg PIXRES_L,
    output reg PIXRES_R,
    output reg STDBY,
    output reg PRECH_COL,
    output reg PGA_RES,
    output reg CK_PH1,
    output reg SAMP_S,
    output reg SAMP_R,
    output reg READ_R,
    output reg READ_S,
    output reg MUX_START,
    output reg CP_COLMUX_IN,
	 output reg DRAIN,
	 output reg PIXGLOB_RES,
    input CLK100MHz,
    input trigger,
	 output reg trigger_ack,
    input [6:0] T1, //times in units of clk100mhz periods (10ns), using ports instead of parameters so no need to resynthesize for optimization 
    input [9:0] T2,
    input [5:0] T3,
    input [9:0] T4,
    input [7:0] T5L,
	 input [7:0] T5R,
    input [4:0] T6,
    input [4:0] T7,
    input [5:0] T8,
    input [6:0] T9,
    input [3:0] T10,
	 input RESET,
	 input ADC_CLKOUT, //3x faster than ADC_PIXCLK, data read clock generated by ADC
	 output ADC_DATA_VALID, //ADC producing valid data, true Tlat3 ADC_CLKOUT cycles after data is collected
	 output ADC_PIXCLK //20MHz PIXCLK to ADCs, trigger synchronized to PIXCLK
    );
	
	parameter Tpix = 10; //time to read 1 pixel, in CLK100MHz periods
	parameter NCOL = 48; //number of columns
	parameter NROW = 176; //number of rows
	parameter Tlat3 = 24;  //number of ADC_CLKOUT cycles before data from a read is output
	
	parameter SM_idle = 1;
	parameter SM_error = 0;
	parameter SM_starting = 2;
	parameter SM_first_signal = 4;
	parameter SM_first_reset = 8;
	parameter SM_left_signal = 16;
	parameter SM_left_reset = 32;
	parameter SM_right_signal = 64;
	parameter SM_right_reset = 128;
	parameter SM_last = 256;
	parameter SM_pixReset = 512;
	
	reg [9:0] timing_SM;
	reg [14:0] counter;
	
	initial timing_SM = SM_idle;
	
	// DCM_SP: Digital Clock Manager
   //         Spartan-6
   // Xilinx HDL Language Template, version 14.7
	wire CLK0;

   DCM_SP #(
      .CLKDV_DIVIDE(Tpix/2),                   // CLKDV divide value
                                            // (1.5,2,2.5,3,3.5,4,4.5,5,5.5,6,6.5,7,7.5,8,9,10,11,12,13,14,15,16).
      .CLKFX_DIVIDE(Tpix/2),                     // Divide value on CLKFX outputs - D - (1-32)
      .CLKFX_MULTIPLY(3),                   // Multiply value on CLKFX outputs - M - (2-32)
      .CLKIN_DIVIDE_BY_2("FALSE"),          // CLKIN divide by two (TRUE/FALSE)
      .CLKIN_PERIOD(10.0),                  // Input clock period specified in nS
      .CLKOUT_PHASE_SHIFT("NONE"),          // Output phase shift (NONE, FIXED, VARIABLE)
      .CLK_FEEDBACK("1X"),                  // Feedback source (NONE, 1X, 2X)
      .DESKEW_ADJUST("SYSTEM_SYNCHRONOUS"), // SYSTEM_SYNCHRNOUS or SOURCE_SYNCHRONOUS
      .DFS_FREQUENCY_MODE("LOW"),           // Unsupported - Do not change value
      .DLL_FREQUENCY_MODE("LOW"),           // Unsupported - Do not change value
      .DSS_MODE("NONE"),                    // Unsupported - Do not change value
      .DUTY_CYCLE_CORRECTION("TRUE"),       // Unsupported - Do not change value
      .FACTORY_JF(16'hc080),                // Unsupported - Do not change value
      .PHASE_SHIFT(0),                      // Amount of fixed phase shift (-255 to 255)
      .STARTUP_WAIT("FALSE")                // Delay config DONE until DCM_SP LOCKED (TRUE/FALSE)
   )
   DCM_SP_ADC(
      .CLK0(CLK0),         // 1-bit output: 0 degree clock output
      //.CLK180(CLK180),     // 1-bit output: 180 degree clock output
      //.CLK270(CLK270),     // 1-bit output: 270 degree clock output
      //.CLK2X(CLK2X),       // 1-bit output: 2X clock frequency clock output
      //.CLK2X180(CLK2X180), // 1-bit output: 2X clock frequency, 180 degree clock output
      //.CLK90(CLK90),       // 1-bit output: 90 degree clock output
      .CLKDV(ADC_PIXCLK),       // 1-bit output: Divided clock output
      //.CLKFX(ADC_INCLK),       // 1-bit output: Digital Frequency Synthesizer output (DFS)
      //.CLKFX180(CLKFX180), // 1-bit output: 180 degree CLKFX output
      //.LOCKED(LOCKED),     // 1-bit output: DCM_SP Lock Output
      //.PSDONE(PSDONE),     // 1-bit output: Phase shift done output
      //.STATUS(STATUS),     // 8-bit output: DCM_SP status output
      .CLKFB(CLK0),       // 1-bit input: Clock feedback input
      .CLKIN(CLK100MHz),       // 1-bit input: Clock input
      .DSSEN(1'b0),       // 1-bit input: Unsupported, specify to GND.
      //.PSCLK(PSCLK),       // 1-bit input: Phase shift clock input
      //.PSEN(PSEN),         // 1-bit input: Phase shift enable
      //.PSINCDEC(PSINCDEC), // 1-bit input: Phase shift increment/decrement input
      .RST(1'b0)            // 1-bit input: Active high reset input
   );

   // End of DCM_SP_inst instantiation
	
	reg ADC_read;
	reg [Tlat3:0] ADC_delay;
	initial ADC_delay = 0;
	reg trigger_sync; //trigger synchronized with ADC_PIXCLK used to signal FSM to start
	initial trigger_sync = 0;
	always@(posedge ADC_CLKOUT)	ADC_delay <= { ADC_read, ADC_delay[Tlat3:1]}; 
	assign ADC_DATA_VALID = ADC_delay[0];
	always@(posedge ADC_PIXCLK) trigger_sync <= trigger;
	
	always @(negedge CLK100MHz) begin
		if (RESET) begin
			timing_SM <= SM_idle;
			ROWADD <= 0;
			COL_L_EN <= 1;
			PIXRES_L <= 1;
			PIXRES_R <= 1;
			STDBY <= 0;
			PRECH_COL <= 0;
			PGA_RES <= 1;
			CK_PH1 <= 0;
			SAMP_S <= 0;
			SAMP_R <= 0;
			READ_R <= 0;
			READ_S <= 0;
			MUX_START <= 1;
			CP_COLMUX_IN <= 1;
			DRAIN <= 0;
			PIXGLOB_RES <= 1;
			counter <= 0;
			trigger_ack <= 0;
			ADC_read <= 0;
		end else begin
			case (timing_SM)  //see timing diagram for state waveforms, this just makes them.
				SM_idle: begin
					ROWADD <= 0;
					COL_L_EN <= 1;
					PIXRES_L <= 0;
					PIXRES_R <= 0;
					STDBY <= 1;
					PRECH_COL <= 0;
					PGA_RES <= 0;
					CK_PH1 <= 0;
					SAMP_S <= 0;
					SAMP_R <= 0;
					READ_R <= 1;
					READ_S <= 0;
					MUX_START <= 1;
					CP_COLMUX_IN <= 1;
					DRAIN <= 0;
					PIXGLOB_RES <= 0;
					trigger_ack <= 0;
					ADC_read <= 0;
					if (trigger_sync) begin 
						timing_SM <= SM_starting;
						/*case(T2%5)
							1:counter <= T2 + 2;  
							2:counter <= T2 + 1;
							3:counter <= T2 + 0;
							4:counter <= T2 + 4;
							default: counter <= T2 + 3;
						endcase*/
						counter <= T2 + Tpix - 2 - (T2 % (Tpix/2)); //the extra time is to make ADC_PIXCLK properly match the read cycle
					end
				end
				SM_starting: begin
					ROWADD <= 0;
					COL_L_EN <= 1;
					PIXRES_L <= 0;
					PIXRES_R <= 0;
					STDBY <= (T2 - 1) < counter;
					PRECH_COL <= 0;
					PGA_RES <= 0;
					CK_PH1 <= 0;
					SAMP_S <= 0;
					SAMP_R <= 0;
					READ_R <= 1;
					READ_S <= 0;
					MUX_START <= 1;
					CP_COLMUX_IN <= 1;
					DRAIN <= 0;
					PIXGLOB_RES <= 0;
					trigger_ack <= 1;
					ADC_read <= 0;
					if (counter == 0) timing_SM <= SM_first_signal;
					else counter <= counter - 1;
				end
				SM_first_signal: begin
					ROWADD <= 0;
					COL_L_EN <= 1;
					PIXRES_L <= 0;
					PIXRES_R <= 0;
					STDBY <= 0;
					PRECH_COL <= counter <= T3;
					PGA_RES <= counter <= T4;
					CK_PH1 <= (T4 < counter) & ((Tpix*NCOL/2 - counter + ((counter - T4) % T5L)) >= T5L) & (((counter - T4) % T5L) < (T5L/2));
					SAMP_S <= T6 <= counter;
					SAMP_R <= 0;
					READ_R <= 1;
					READ_S <= 0;
					MUX_START <= 1;
					CP_COLMUX_IN <= 1;
					DRAIN <= 1;
					PIXGLOB_RES <= 0;
					trigger_ack <= 1;
					ADC_read <= 0;
					if (counter >= Tpix*NCOL/2) begin
						timing_SM <= SM_first_reset;
						counter <= 1;
					end else counter <= counter + 1;
				end
				SM_first_reset: begin
					ROWADD <= 0;
					COL_L_EN <= 1;
					PIXRES_L <= counter <= T1;
					PIXRES_R <= 0;
					STDBY <= 0;
					PRECH_COL <= 0;
					PGA_RES <= counter <= T4;
					CK_PH1 <= (T4 < counter) & ((Tpix*NCOL/2 - counter + ((counter - T4) % T5L)) >= T5L) & (((counter - T4) % T5L) < (T5L/2));
					SAMP_S <= 0;
					SAMP_R <= T6 <= counter;
					READ_R <= 1;
					READ_S <= 0;
					MUX_START <= 1;
					CP_COLMUX_IN <= 1;
					DRAIN <= 1;
					PIXGLOB_RES <= 0;
					trigger_ack <= 1;
					ADC_read <= 0;
					if (counter >= Tpix*NCOL/2) begin
						timing_SM <= SM_right_signal;
						counter <= 1;
					end else counter <= counter + 1;
				end
				SM_right_signal: begin
					ROWADD <= ROWADD;
					COL_L_EN <= 0;
					PIXRES_L <= 0;
					PIXRES_R <= 0;
					STDBY <= 0;
					PRECH_COL <= counter <= T3;
					PGA_RES <= counter <= T4;
					CK_PH1 <= (T4 < counter) & ((Tpix*NCOL/2 - counter + ((counter - T4) % T5R)) >= T5R) & (((counter - T4) % T5R) < (T5R/2));
					SAMP_S <= T6 <= counter;
					SAMP_R <= 0;
					READ_R <= (counter % Tpix) < T8;
					READ_S <= ((T7 + T8) <= (counter % Tpix)) & ((counter % Tpix) < (T8 + T7 + T8));
					MUX_START <= counter <= T9;
					CP_COLMUX_IN <= (((T7 + T8 + T8 + T10) % Tpix) <= (counter % Tpix)) & ((counter % Tpix) < ((T7 + T8 + T8 + T10 + 4) % Tpix));
					DRAIN <= 1;
					PIXGLOB_RES <= 0;
					trigger_ack <= 1;
					ADC_read <= 1;
					if (counter >= Tpix*NCOL/2) begin
						timing_SM <= SM_right_reset;
						counter <= 1;
					end else counter <= counter + 1;
				end
				SM_right_reset: begin
					ROWADD <= ROWADD;
					COL_L_EN <= 0;
					PIXRES_L <= 0;
					PIXRES_R <= counter <= T1;
					STDBY <= 0;
					PRECH_COL <= 0;
					PGA_RES <= counter <= T4;
					CK_PH1 <= (T4 < counter) & ((Tpix*NCOL/2 - counter + ((counter - T4) % T5R)) >= T5R) & (((counter - T4) % T5R) < (T5R/2));
					SAMP_S <= 0;
					SAMP_R <= T6 < counter;
					READ_R <= (counter % Tpix) < T8;
					READ_S <= ((T7 + T8) <= (counter % Tpix)) & ((counter % Tpix) < (T8 + T7 + T8));
					MUX_START <= 0;
					CP_COLMUX_IN <= (((T7 + T8 + T8 + T10) % Tpix) <= (counter % Tpix)) & ((counter % Tpix) < ((T7 + T8 + T8 + T10 + 4) % Tpix));
					DRAIN <= 1;
					PIXGLOB_RES <= 0;
					trigger_ack <= 1;
					ADC_read <= 1;
					if (counter >= Tpix*NCOL/2) begin
						timing_SM <= (ROWADD == NROW - 1)?SM_last:SM_left_signal;
						counter <= 1;
					end else counter <= counter + 1;
				end
				SM_left_signal: begin
					if (counter == 1) ROWADD <= ROWADD + 1;
					else ROWADD <= ROWADD;
					COL_L_EN <= 1;
					PIXRES_L <= 0;
					PIXRES_R <= 0;
					STDBY <= 0;
					PRECH_COL <= counter <= T3;
					PGA_RES <= counter <= T4;
					CK_PH1 <= (T4 < counter) & ((Tpix*NCOL/2 - counter + ((counter - T4) % T5L)) >= T5L) & (((counter - T4) % T5L) < (T5L/2));
					SAMP_S <= T6 < counter;
					SAMP_R <= 0;
					READ_R <= (counter % Tpix) < T8;
					READ_S <= ((T7 + T8) <= (counter % Tpix)) & ((counter % Tpix) < (T8 + T7 + T8));
					MUX_START <= counter <= T9;
					CP_COLMUX_IN <= (((T7 + T8 + T8 + T10) % Tpix) <= (counter % Tpix)) & ((counter % Tpix) < ((T7 + T8 + T8 + T10 + 4) % Tpix));
					DRAIN <= 1;
					PIXGLOB_RES <= 0;
					trigger_ack <= 1;
					ADC_read <= 1;
					if (counter >= Tpix*NCOL/2) begin
						timing_SM <= SM_left_reset;
						counter <= 1;
					end else counter <= counter + 1;
				end
				SM_left_reset: begin
					ROWADD <= ROWADD;
					COL_L_EN <= 1;
					PIXRES_L <= counter <= T1;
					PIXRES_R <= 0;
					STDBY <= 0;
					PRECH_COL <= 0;
					PGA_RES <= counter <= T4;
					CK_PH1 <= (T4 < counter) & ((Tpix*NCOL/2 - counter + ((counter - T4) % T5L)) >= T5L) & (((counter - T4) % T5L) < (T5L/2));
					SAMP_S <= 0;
					SAMP_R <= T6 < counter;
					READ_R <= (counter % Tpix) < T8;
					READ_S <= ((T7 + T8) <= (counter % Tpix)) & ((counter % Tpix) < (T8 + T7 + T8));
					MUX_START <= 0;
					CP_COLMUX_IN <= (((T7 + T8 + T8 + T10) % Tpix) <= (counter % Tpix)) & ((counter % Tpix) < ((T7 + T8 + T8 + T10 + 4) % Tpix));
					DRAIN <= 1;
					PIXGLOB_RES <= 0;
					trigger_ack <= 1;
					ADC_read <= 1;
					if (counter >= Tpix*NCOL/2) begin
						timing_SM <= SM_right_signal;
						counter <= 1;
					end else counter <= counter + 1;
				end
				SM_last: begin
					ROWADD <= NROW;
					COL_L_EN <= 1;
					PIXRES_L <= 0;
					PIXRES_R <= 0;
					STDBY <= 0;
					PRECH_COL <= 0;
					PGA_RES <= 0;
					CK_PH1 <= 0;
					SAMP_S <= 0;
					SAMP_R <= 0;
					READ_R <= (counter % Tpix) < T8;
					READ_S <= ((T7 + T8) < (counter % Tpix)) & ((counter % Tpix) < (T8 + T7 + T8));
					MUX_START <= counter <= T9;
					CP_COLMUX_IN <= (((T7 + T8 + T8 + T10) % Tpix) < (counter % Tpix)) & ((counter % Tpix) < ((T7 + T8 + T8 + T10 + 4) % Tpix));
					DRAIN <= 1;
					PIXGLOB_RES <= 0;
					trigger_ack <= 1;
					ADC_read <= 1;
					if (counter >= Tpix*NCOL/2) begin
						timing_SM <= SM_pixReset;
						counter <= 1;
					end else counter <= counter + 1;
				end
				SM_pixReset: begin
					ROWADD <= NROW;
					COL_L_EN <= 1;
					PIXRES_L <= 0;
					PIXRES_R <= 0;
					STDBY <= 1;
					PRECH_COL <= 0;
					PGA_RES <= 0;
					CK_PH1 <= 0;
					SAMP_S <= 0;
					SAMP_R <= 0;
					READ_R <= 1;
					READ_S <= 0;
					MUX_START <= 1;
					CP_COLMUX_IN <= 1;
					DRAIN <= 1;
					PIXGLOB_RES <= 1;
					trigger_ack <= 1;
					ADC_read <= 0;
					if (counter == Tpix*NCOL/2) begin
						timing_SM <= SM_idle;
						counter <= 0;
					end else counter <= counter + 1;
				end
			endcase
		end
	end
	
endmodule
